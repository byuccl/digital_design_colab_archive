module add_8(
  input logic cin,
  input logic [7:0] a, b,
  output logic [7:0] s,
  output logic co 
  );
  //Instantiate 8 instances of full_adder
  //Have cin be the first carry in and co be the last carry out
  
 endmodule
