module mod_counter#(
  //Add the parameter
)(
  //Add the Inputs exactly as listed
);
  //Code
endmodule
