module seven_segment_top (
  input logic [3:0] sw,
  input logic btnc,
  output logic [7:0] segment,
  output logic [3:0] anode
);

  //Top module for seven_segment
  
endmodule
