module stopwatch(
  //Signals
);
  //Code
endmodule
