module stopwatch_top (
  //Signals
);
endmodule
