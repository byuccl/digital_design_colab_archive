module function1 (
 output logic [15:0] led,
 input logic  btnd,
 input logic [15:0] sw
);
    
// Code goes here

endmodule // behavLoadableReg
