module full_add(
  input logic a, b, cin,
  output logic s, co
  );
  //A, B and the cin should be added together. s is the result and co signifies carry over.
  endmodule
