module seven_segment(
  input logic [3:0] data,
  output logic [6:0] segment
);
  //Data should be converted into seven segment signals
  
endmodule
